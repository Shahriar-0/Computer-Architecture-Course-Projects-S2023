module RegID_EX();

endmodule