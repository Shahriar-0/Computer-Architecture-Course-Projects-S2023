module ForwardingUnit();

endmodule