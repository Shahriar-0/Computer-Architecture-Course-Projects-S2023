module RegMEM_WB();

endmodule