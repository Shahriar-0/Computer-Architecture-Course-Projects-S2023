module RegIF_ID();

endmodule