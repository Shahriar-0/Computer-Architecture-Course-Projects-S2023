module ALU_Controller(op, func, aluOp);

    input [1:0] op;
    input [5:0] func;

    output reg [2:0] aluOp;
    
endmodule
