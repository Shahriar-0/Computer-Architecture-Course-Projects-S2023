timescale 1ns / 1ns

module tb();

    intelligent_rat rat;
    initial begin
        // sth
    end

endmodule