module InstructionMemory (pc, instruction);
    input [31:0] pc;
    output [31:0] instruction;

    
endmodule
