module BranchController (branch, zero, pcSrc);
    input branch, zero;
    output reg pcSrc;
    reg pcSrc;

    
endmodule