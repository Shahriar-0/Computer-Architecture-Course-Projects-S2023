`timescale 1ns/1ns

module datapath(input CLK,RST,init_x,init_y,ld_x,ld_y,ld_count,init_count,en_count,list_push,list_read,
    init_read_ptr,stack_dir_push,stack_dir_pop,r_update,output_x,output finish,empty_stack,list_empty,Co);



endmodule