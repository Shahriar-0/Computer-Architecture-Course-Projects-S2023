module RegEX_MEM();

endmodule