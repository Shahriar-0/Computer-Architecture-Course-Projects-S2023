module RISC_V_Controller(); 

endmodule