module HazardUnit();

endmodule